module hub75_driver (
    input wire clk_in,

    output wire R0,
    output wire R1,
    output wire G0,
    output wire G1,
    output wire B0,
    output wire B1,

    output wire A,
    output wire B,
    output wire C,
    output wire D,
    output wire E,

    output wire CLK,
    output wire STB,
    output wire OE
);
    // TODO: Literally everything!
endmodule
