module divider (
	input [31:0] dividend,
	input [31:0] divisor,
	input wire signed,
	output [31:0] quotient,
	output [31:0] remainder,
);
	
endmodule